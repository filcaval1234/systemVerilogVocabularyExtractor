`include "tb_diff.sv"
